library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;
use work.functions.all;

entity demodulate is
generic
(
	GAIN: natural:= 0
	);
port
(
	clock: in std_logic;
	reset: in std_logic;
	real_in : in std_logic_vector (31 downto 0);
    imag_in : in std_logic_vector (31 downto 0);
    real_empty : in std_logic;
    imag_empty : in std_logic;
    out_full : in std_logic;
    real_rd_en : out std_logic;
    imag_rd_en : out std_logic;
    dout : out std_logic_vector (31 downto 0);
    out_wr_en : out std_logic
    );
end entity;

type states is(init, read, divide, write);
signal state,next_state:states:=init;
signal real_prev,real_prev_c,imag_prev,imag_prev_c: stdlogic_vector(31 downto 0);
signal divisor,divisor_c,dividend,dividend_c,quotient,quotient_c: signed(31 downto 0);
signal quad_a,quad_a_c,quad_b,quad_b_c:integer:=0;
signal a,a_c,b,b_c,q,q_c,y,y_c:signed(31 downto 0);
 demod_process : process (state, real_prev, imag_prev, dividend, divisor, quotient, quad_a, quad_b, a, b, q, y, real_in, imag_in, real_empty, imag_empty, out_full)
        variable r, i : signed (31 downto 0) := (others => '0');
        variable dividend_v, divisor_v : signed (31 downto 0) := (others => '0');
        variable p : integer := 0;
        variable sign : std_logic := '0';
		variable angle : signed (31 downto 0) := (others => '0');
		begin
	    next_state <= state;
        real_prev_c <= real_prev;
        imag_prev_c <= imag_prev;
        dividend_c <= dividend;
        divisor_c <= divisor;
        quotient_c <= quotient;
        quad_a_c <= quad_a;
        quad_b_c <= quad_b;
        a_c <= a;
        b_c <= b;
        q_c <= q;
        y_c <= y;

        real_rd_en <= '0';
        imag_rd_en <= '0';
        out_wr_en <= '0';
        dout <= (others => '0');

        dividend_v := (others => '0');
        divisor_v := (others => '0');
        angle := (others => '0');

        case (state) is
            when init =>
                if (real_empty = '0' and imag_empty = '0') then
                    real_prev_c <= (others => '0');
                    imag_prev_c <= (others => '0');
                    dividend_c <= (others => '0');
                    divisor_c <= (others => '0');
                    quotient_c <= (others => '0');
                    a_c <= (others => '0');
                    b_c <= (others => '0');
                    q_c <= (others => '0');
                    quad_a_c <= 0;
                    quad_b_c <= 0; 
                    y_c <= (others => '0');
                    next_state <= read;
                end if;

               when read =>
                if (real_empty = '0') then
                    dividend_c <= (others => '0');
                    divisor_c <= (others => '0');
                    quotient_c <= (others => '0');
                    a_c <= (others => '0');
                    b_c <= (others => '0');
                    q_c <= (others => '0');
                    quad_a_c <= 0;
                    quad_b_c <= 0; 
                    y_c <= (others => '0');

                    real_rd_en <= '1';
                    imag_rd_en <= '1';

                    r := DEQUANTIZE(signed(real_in) * signed(real_prev)) - DEQUANTIZE(-signed(imag_prev) * signed(imag_in));
                    i := DEQUANTIZE(signed(imag_in) * signed(real_prev)) + DEQUANTIZE(-signed(imag_prev) * signed(real_in));
                    y_c <= i;
                    i := abs(i) + 1;

                    real_prev_c <= real_in;
                    imag_prev_c <= imag_in;

                    if (r >= 0) then
                        --angle = QUAD1 - DEQUANTIZE(QUAD1 * DIV(QUANTIZE(r - i), r + i))
                        quad_a_c <= QUAD1;
                        quad_b_c <= QUAD1;
                        dividend_v := QUANTIZE(r - i);
                        divisor_v := r + i;
                    else
                        --angle = QUAD3 - DEQUANTIZE(QUAD3 * DIV(QUANTIZE(r + i), i - r))
                        quad_a_c <= QUAD3; 
                        quad_b_c <= QUAD1;
                        dividend_v := QUANTIZE(r + i);
                        divisor_v := i - r;
                    end if;

                    dividend_c <= dividend_v;
                    divisor_c <= divisor_v;
                    a_c <= abs(dividend_v);
                    b_c <= abs(divisor_v);

                    next_state <= divide;
                end if;

            when divide =>
                if (b = 1) then
                    q_c <= a;
                    a_c <= (others => '0'); 
                end if;

                if (a >= b) then
                    p := GET_MSB(signed(a)) - GET_MSB(signed(b));
                    if ((b sll p) > a) then
                        p := p - 1;
                    end if;
                    q_c <= q + (to_signed(1, WORD) sll p);
                    a_c <= a - (b sll p);
                else
                    quotient_c <= q; 
                    sign := dividend(31) xor divisor(31);
                    if (sign = '1') then
                        quotient_c <= -q; 
                    end if;
                    next_state <= write;
                end if;

            when write =>
                if (demod_full = '0') then
                    angle := quad_a - DEQUANTIZE(quad_b * quotient);
                    if (y < 0) then
                        angle := -angle;
                    end if;
                    dout <= std_logic_vector(DEQUANTIZE(GAIN * angle));
                    out_wr_en <= '1';
                    next_state <= read;
                end if;

            when others =>
                next_state <= init;

        end case;
    end process;

    clock_process : process (clock, reset)
    begin 
        if (reset = '1') then
            state <= init;
            real_prev <= (others => '0'); 
            imag_prev <= (others => '0'); 
            dividend <= (others => '0');  
            divisor <= (others => '0');  
            quotient <= (others => '0');  
            quad_a <= 0; 
            quad_b <= 0; 
            a <= (others => '0'); 
            b <= (others => '0'); 
            q <= (others => '0'); 
            y <= (others => '0'); 
        elsif (rising_edge(clock)) then
            state <= next_state;
            real_prev <= real_prev_c;
            imag_prev <= imag_prev_c;
            dividend <= dividend_c;
            divisor <= divisor_c;
            quotient <= quotient_c;
            quad_a <= quad_a_c;
            quad_b <= quad_b_c;
            a <= a_c;
            b <= b_c;
            q <= q_c;
            y <= y_c;
        end if;
    end process;

end architecture;
